`timescale 1ns / 1ps

module positadd_tb;
    parameter N = 32;
    parameter es = 3;

    reg [N-1:0] in1, in2;
    reg start;
    wire [N-1:0] out;
    wire done;
    reg clk;

    // Instantiate the Unit Under Test (UUT)
    positadd_4_es3 uut (
        .clk(clk),
        .in1(in1),
        .in2(in2),
        .start(start),
        .result(out),
        .inf(inf),
        .zero(zero),
        .done(done)
    );

	initial
    begin
		// Initialize Inputs
		in1 = 0;
		in2 = 0;
		clk = 0;
		start = 1;

        in1 = 32'b00101100011010110100010000111011;
        in2 = 32'b11001011011001101111101111111001;
        // 11001101000000111001101000010000

        // 1 01 100 10111111000110010111110000


	end

    always #5
    begin
        clk = ~clk;
    end
endmodule
