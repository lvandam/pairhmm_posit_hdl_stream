// Right shift unit
module DSR_right_N_S(a, b, c);
    parameter N = 16;
    parameter S = 4;
    
    input [N-1:0] a;
    input [S-1:0] b;
    output [N-1:0] c;

    wire [N-1:0] tmp [S-1:0];
    assign tmp[0] = b[0] ? (a >> 7'd1) : a;

    genvar i;
    generate
    	for (i = 1; i < S; i = i + 1)
        begin: loop_blk
    		assign tmp[i] = b[i] ? (tmp[i-1] >> 2**i) : tmp[i-1];
    	end
    endgenerate

    assign c = tmp[S-1];

endmodule
