module add_mantovf (a, mant_ovf, c);
    parameter N = 10;
    input [N:0] a;
    input mant_ovf;
    output [N:0] c;

    assign c = a + mant_ovf;
endmodule
